BSV1    T�k��1  NESS����TIME   (   +}  CPUR   W����  PPUR4   �� �    ")60!' ' 0' 0' 6t�t�    APURH   �j�� �	 0  �   ^     jJ     $     
    ��    �    CTRL   ��������    MAPR    LRAM    � p   �                                                            ����                                  rp�����                                                         ��x���                   ���       [�"                             i      �             0                                                   ������������������������������������������������������������������������������������������������������������������������������������������=��=��o� O ��W��#X�  p�! x�" p�# x�$ p�% x�& p�' x�   ��C���C��qC��pC��sC��rC���Cø�C��qC��pC��sC��rC˸�Cڸ�C��qC��pC��sC��rC��sC��rC���C���C��qC��pC��sC��rC���C���C��qC��pC���!���a���!���a���!���a���C���C��qC��pC��sC��rC���C���C��qC��pC��sC��rC�x�!�x�a���!���a���!���a�  ' z                                                    � '� '� '� '� '�T'�                                                                   �            p�         ��                                                                     p�  �                 �xx� x                        ��                          �                                                              �         					             r�~����������Ƹ���������                                                                                                         ��                                                   �                                                                     TTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTT                                                                                                         �                                                          TTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTT         NTT                                                XH8��(@Xp���$����X`hpx����     �( ����            � $�    &  $���                    B   p   O   F Y          ""                	   	                          hn�c��  r  	    @ 0p    k                                            	     �SPRT   �#X�  p�! x�" p�# x�$ p�% x�& p�' x�   ��C���C��qC��pC��sC��rC���Cø�C��qC��pC��sC��rC˸�Cڸ�C��qC��pC��sC��rC��sC��rC���C���C��qC��pC��sC��rC���C���C��qC��pC���!���a���!���a���!���a���C���C��qC��pC��sC��rC���C���C��qC��pC��sC��rC�x�!�x�a���!���a���!���a�NTAB   $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$
$$$$$$$$$$ $$$$$$$$$$$$ $$.) $$$$($$$$ $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$6767$$$$$$$$$$$$$$$$$$$$$$$$$$$5%%%%8$$$$$$$$$$$$$$$$$$$$$$$$$$9:;:;<$$$$$$$$$$$$$$$$$$$����$$$$$$$$$$$$$$$$$$$$$$$$$$$$����$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$��$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$��$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$`abc$$$$$$$$$$$$$$$$$$$$$$$$$$$$defg$$$$$$$$$$$$$$$$$$$$$$$$$$$$hi&j$$$$$$��$$$$$$$$$$$$$$$$$$$$hi&j$$$$$$��$$$$$$$$$$$$$$$$$$$$hi&j$$��$$��$$$$$$$$$$$$$$$$$$$$hi&j$$��$$��$$$$$$$$$$$$$$$$$$$$hi&j$$��$$������$$$$$$$$$$$$$$$$hi&j$$��$$����������������������������������������������������������������������������������������������������������������������������������������ꪪ�����      

                           PPPPPTTU$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$67$$$$$$$$$$$$$$$$$$$$$$$$$$$$$5%%8$$$$$$$67$$$$$$$$$$$$$$$$$$$9:;<$$$$$$5%%8$$$$$$$$$$$$$$$$$$$$$$$$$$$$9:;<$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$��$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$��$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$`abc$$$$$$$$$$$$$$$$$$$$$$$$$$$$defg$$$$$$$$$$��$$$$$$$$$$��$$$$hi&j$$$$$$$$$$��$$$$$$$$$$��$$$$hi&j$$$$$$`abc��$$����$$$$��$$$$hi&j$$$$$$defg��$$����$$$$��$$$$hi&j����$$hi&j��$$������$$��$$$$hi&j����$$hi&j��$$������$$��$$$$hi&j��������������������������������������������������������������������������������������������������������������������������������         �    �� 
                            UPTTUTPPSRAM    ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������gend                                                                                                                                                                                                                                                                                                                                                                    