BSV1    D��d�1  NESS����TIME      �M  CPUR   W����  PPUR4   �� �     ")60! ' 0' 0' 6n�n�    APURH   �j�� |	 X0  �   [      y                sQ{    �    CTRL   ��������    MAPR    LRAM   � J   ?@  @                                                                  �                                        JPPPP                   �                                            �n                       ��N�       �                                                                                                      �������������������������������������������������������������������������������������������������������������������������������������������==��=��o� O ��W��#X��@J��@R��@J��@R�A@J�2@R�C@J�B@R�   �   �   ��A�iA��A�jA��A��A�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ��A�iA��A�jA��A��A�   �   �   �   �   �   �   �   �   �   �   �   ��A�iA��A�jA��A��A�   �   �   �   �   �      '                                                                                                                                                 �            J         �n                                                                     �                    $T                           �,                           �                                                              �                         M�W�����                                                                                                                                                                                                                                                            TTTTTTTTTTTTTTT TTTTTTTTTTTTTTT                                                                        a              aa              aa            a aa           aa aa          aaa aa         aaaa aa        TTTTT TT        TTTTT TT            aaaaaaaTT                                     �          XH8�����(@Xh$x|�����(08@HP   0  0�``               �� $�       
���                     2  J    M  /Y          ""                 
                              ���Yu  $        0!    X                                          		    �SPRT   �#X��@J��@R��@J��@R�A@J�2@R�C@J�B@R�   �   �   ��A�iA��A�jA��A��A�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ��A�iA��A�jA��A��A�   �   �   �   �   �   �   �   �   �   �   �   ��A�iA��A�jA��A��A�   �   �   �   �   �   NTAB   $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$
$$$$$$$$$$ $$$$$$$$$$$$$$.)$$$$($$$$		$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$6767$$$$$$$$$$$$$$$$$$$$$$$$$$$5%%%%8$$$$$$$$$$$$$$$$$$$$$$$$$$9:;:;<$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$������$$$$$$$$$$$$$$$$$$$$$$$$$$GGGGGG$$$$$$$$$$$$$$$$$$$$$$$$$$G'GG'G$$$$$$$$$$$$$$$$$$$$$$$$$$G'GG'G$$$$$$$$$$$$$$$$$$$$$$$$����������$$$$$$$$$$$$$$$$��$$$$GGGGGGGGGG$$$$$$$$$$$$$$$$��$$$$GGGG��GGGG$$$$$$$$$$$$��$$��$$$$GGGG''GGGG$$$$$$$$$$$$��$$��$$$$GGGG''GGGG$$$$$$$$$$$$��$$����$$GGGG''GGGG$$$$$$$$$$$$��$$����$$������������������������������$$������������������������������$$������������������������������$$������������������������������$$��ꪪ�����      

              DU      UU     UUQPPTT$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$67$$$$$$$$$$$$$$$$$$$$$$$$$$$$$5%%8$$$$$$$$$$$$$$$$$$$$$$$$$$$$9:;<$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$��$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$��$$$$$$$$$$$$$$$$$$$$$$$$$$$$����$$$$$$$$$$$$$$$$$$$$$$$$$$$$����$$$$$$$$$$$$$$$$$$$$$$$$$$$$����$$$$$$$$$$$$$$$$$$$$$$$$$$$$����$$$$$$$$$$$$$$$$$$$$$$$$��$$����$$$$$$$$$$$$$$$$$$$$$$$$��$$����$$$$$$$$$$$$$$$$$$$$$$����$$����$$$$$$$$$$$$$$$$$$$$$$����$$����$$$$$$$$$$$$$$$$$$$$������$$����$$$$$$$$$$$$$$$$$$$$������$$����$$$$$$$$$$$$$$$$����������$$����$$$$$$$$$$$$$$$$����������$$����$$$$$$$$$$$$$$$$����������$$����$$$$$$$$$$$$$$$$����������$$����$$$$$$$$$$$$$$$$����������$$����$$$$$$$$$$$$$$$$����������$$����$$$$$$$$$$$$$$$$         �       
        T      U     TU    UUU        SRAM    ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������gend                                                                                                                                                                                                                                                                                                                                                                                                                                                                